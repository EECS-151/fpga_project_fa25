`timescale 1ns/1ns

module counter_tb();

// TODO: Use the other testbenches and your counter_testbench from Lab 2 as a guide

endmodule